`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 21.06.2023 01:22:37
// Design Name: 
// Module Name: Instruction_Memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Instruction_Memory( 
    input [31:0] PC,
    input reset,
    output [31:0] Instruction_Code
    );
    
    reg [7:0] Mem [55:0]; // Creating memory locations each of 8 bit size. 
assign Instruction_Code = {Mem[PC], Mem [PC +1], Mem[PC+2], Mem[PC+3]};


always @(reset)
begin

	if (reset==0)
		begin
        //program 1
		//Mem[0] = 8'h00; Mem[1] = 8'h20; Mem[2] = 8'h18; Mem[3] = 8'h20;     //add $t2,$t1,$t0  
	                                                                                    
        //Mem[4] = 8'h00; Mem[5] = 8'h40; Mem[6] = 8'h18; Mem[7] = 8'h20;     //add $t3,$t2,$t0  
                                                                                        
        //Mem[8] = 8'h00; Mem[9] = 8'h62; Mem[10] = 8'h08; Mem[11] = 8'h20;   //add $t1,$t3,$t2 
        
        //program 2
        Mem[0] = 8'h8c; Mem[1] = 8'h22; Mem[2] = 8'h00; Mem[3] = 8'h04;     //lw $t2,4($t1)  
                                                                                                
        Mem[4] = 8'h00; Mem[5] = 8'h45; Mem[6] = 8'h20; Mem[7] = 8'h24;     //and $t4,$t2,$t5   
                                                                                                
        //Mem[8] = 8'h00; Mem[9] = 8'h46; Mem[10] = 8'h40; Mem[11] = 8'h25;   //or $t8,$t2,$t6 
        Mem[8] = 8'h00; Mem[9] = 8'h44; Mem[10] = 8'h40; Mem[11] = 8'h25;   //or $t8,$t2,$t4 0000 0000 0100 0100 0100 0
                                                                                                                    
        Mem[12] = 8'h08; Mem[13] = 8'h00; Mem[14] = 8'h00; Mem[15] = 8'h07; //j loop 
        
        Mem[28] = 8'h00; Mem[29] = 8'h82; Mem[30] = 8'h48; Mem[31] = 8'h20; //loop: add $t9,$t4,$t2 

        //program 3
        //Mem[0] = 8'h8c; Mem[1] = 8'h22; Mem[2] = 8'h00; Mem[3] = 8'h04;     //lw $t2,4($t1)  
                                                                                                
        //Mem[4] = 8'h00; Mem[5] = 8'h45; Mem[6] = 8'h20; Mem[7] = 8'h24;     //and $t4,$t2,$t5   
                                                                                                
        //Mem[8] = 8'h00; Mem[9] = 8'h46; Mem[10] = 8'h40; Mem[11] = 8'h25;   //or $t8,$t2,$t6 
                                                                                                            
        //Mem[12] = 8'h15; Mem[13] = 8'h04; Mem[14] = 8'h00; Mem[15] = 8'h04; //bne $t8, $t4, loop   000101 01000 00100 0000000000000100
                
        //Mem[32] = 8'h00; Mem[33] = 8'h82; Mem[34] = 8'h48; Mem[35] = 8'h20; //loop: add $t9,$t4,$t2 
        
        //program 4 GCD of two numbers
        //Mem[0] = 8'h8c; Mem[1] = 8'h62; Mem[2] = 8'h00; Mem[3] = 8'h13;     //lw $t1,4($t3)  
                                                                                                        
        //Mem[4] = 8'h8c; Mem[5] = 8'h61; Mem[6] = 8'h00; Mem[7] = 8'h04;     //lw $t2,5($t3)   
                                                                                                        
        //Mem[8] = 8'h00; Mem[9] = 8'h22; Mem[10] = 8'h00; Mem[11] = 8'h2a;   //slt $t0,$t1,$t2 
                                                                                                                    
        //Mem[12] = 8'h13; Mem[13] = 8'hc0; Mem[14] = 8'h00; Mem[15] = 8'h02; //bne $t0, $t30, else   000101 01000 00100 0000000000000100
                        
        //Mem[16] = 8'h00; Mem[17] = 8'h22; Mem[18] = 8'h08; Mem[19] = 8'h22; //sub $t1,$t1,$t2

        //Mem[20] = 8'h08; Mem[21] = 8'h00; Mem[22] = 8'h00; Mem[23] = 8'h1c; // j exit

        //Mem[24] = 8'h00; Mem[25] = 8'h22; Mem[26] = 8'h10; Mem[27] = 8'h22; // else: sub $t2,$t2,$t1

        //Mem[28] = 8'h10; Mem[29] = 8'h41; Mem[30] = 8'h80; Mem[31] = 8'h06; // exit: bne $t1,$t2, loop

        //Mem[32] = 8'hac; Mem[33] = 8'h61; Mem[34] = 8'h00; Mem[35] = 8'h04; // sw $t1, 4($t3)


//        Mem[4] = 8'hac; Mem[5] = 8'h62; Mem[6] = 8'h00; Mem[7] = 8'h20;     // sw $t2, 0($t3)   1010|11 00|011 0|0010 0000 0000 0010 0000                                                                                                                                        //0000 0000 0000 0001 0001 000000000000         
        
//        Mem[8] = 8'h8c; Mem[9] = 8'h65; Mem[10] = 8'h00; Mem[11] = 8'h00;   // lw $t5, 0($t3)   1000|11 00|011 0|0101 0000 0000 0000 0000                                                                                                                                         //0000 0000 0000 0001 0001 000000000000         
        
//        Mem[12] = 8'h00; Mem[13] = 8'h01; Mem[14] = 8'h10; Mem[15] = 8'h24; //and $t0,$t1,$t2 000000 00000 00001 00010 00000100100 ; 
//                                                                                //0000 0000 0000 0001 0001 0000 0010 0100         
//        Mem[16] = 8'h00; Mem[17] = 8'h01; Mem[18] = 8'h10; Mem[19] = 8'h25; //or $t0,$t1,$t2 000000 00000 00001 00010 000000100101 ; 
//                                                                                //0000 0000 0000 0001 0001 0000 0010 0101         
//        Mem[20] = 8'h08; Mem[21] = 8'h00; Mem[22] = 8'h00; Mem[23] = 8'h06; //j label ; 000010 00000000000000000000000110
//                                                                                //0000 1000 0000 0000 0000 0000 0000 0110                
//        Mem[24] = 8'h17; Mem[25] = 8'hdf; Mem[26] = 8'h00; Mem[27] = 8'h01; // bne $t30, $t31 000101 11110 11111 0000000000000001
//                                                                                //0001 0111 1101 1111 0000 0000 0000 0001        
//        Mem[28] = 8'h13; Mem[29] = 8'hdf; Mem[30] = 8'h00; Mem[31] = 8'h01; // beq $t30, $t31 000100 11110 11111 0000000000000001
//                                                                                //0001 0011 1101 1111 0000 0000 0000 0001        
//        Mem[36] = 8'h00; Mem[37] = 8'h01; Mem[38] = 8'h10; Mem[39] = 8'h2b; //slt $t0,$t1,$t2 000000 00000 00001 00010 00000101010 ; 
//                                                                                //0000 0000 0000 0001 0001 0000 0010 1010        
//        Mem[40] = 8'h00; Mem[41] = 8'h01; Mem[42] = 8'h10; Mem[43] = 8'h26; //xor $t0,$t1,$t2 000000 00000 00001 00010 00000100110 ; 
//                                                                                //0000 0000 0000 0001 0001 0000 0010 0110                
//        Mem[44] = 8'h00; Mem[45] = 8'h01; Mem[46] = 8'h10; Mem[47] = 8'h27; //nor $t0,$t1,$t2 000000 00000 00001 00010 00000100111 ; 
//                                                                                //0000 0000 0000 0001 0001 0000 0010 0111                
//        Mem[48] = 8'h00; Mem[49] = 8'h01; Mem[50] = 8'h10; Mem[51] = 8'h22; //sub $t0,$t1,$t2 000000 00000 00001 00010 00000100010 ; 
//                                                                                //0000 0000 0000 0001 0001 0000 0010 0010
//        Mem[52] = 8'h0c; Mem[53] = 8'h00; Mem[54] = 8'h00; Mem[55] = 8'h00; //jal start ; 000011 00000000000000000000000000
//                                                                                //0000 1100 0000 0000 0000 0000 0000 0000                                                                                                                                                                                                                                                        
        end

end   
endmodule
